(* regbank_gen *)
module regbank();
endmodule
